// SPDX-License-Identifier: BSD-3-clause
/*
 * Copyright (C) Till Mahlburg, 2023
 *
 * Project    : Memory Tagged SEC-V
 * Author     : Till Mahlburg
 * Purpose    : Memory Tagging function unit for the SEC-V processor.
 *
 * TODO:
 *      - use shift operation to calculate tmem_adr_o
 *
 * History
 *    v1.0        - Initial version
 */

`include "secv_pkg.svh"
import secv_pkg::*;

module mtag #(
    /* size of tags in bit */
    parameter int TLEN = 16,
    /* size of granules in byte */
    parameter int GRANULARITY = 8,
    /* address size in bit */
    parameter int ADR_WIDTH = 8,
    /* tag memory address width in bit */
    parameter int TADR_WIDTH = 16,
    /* tag memory byte selection width */
    parameter int TSEL_WIDTH = TLEN / 8
) (
    input funit_in_t fu_i,
    output funit_out_t fu_o,

    /* tag memory */
    output logic                    tmem_cyc_o,
    output logic                    tmem_stb_o,
    output logic [TSEL_WIDTH-1 : 0] tmem_sel_o,
    output logic [TADR_WIDTH-1 : 0] tmem_adr_o,
    output logic                    tmem_we_o,
    output logic [TLEN-1 : 0]       tmem_dat_o,
    input  logic                    tmem_ack_i
);
    logic [ADR_WIDTH-1 : 0] mem_adr;
    assign mem_adr = ADR_WIDTH'(fu_i.src1);

    // decode encoded tag
    logic [TLEN-1 : 0] enc_tag;
    assign enc_tag = fu_i.src1[XLEN-1 : XLEN-TLEN];

    // decode tag from rs2
    logic [TLEN-1 : 0] r_tag;
    assign r_tag = TLEN'(fu_i.src2);

    logic err;

    always_comb begin
        err = 'b0;

        tmem_cyc_o = 'b0;
        tmem_stb_o = 'b0;
        tmem_sel_o = 'b0;
        tmem_adr_o = 'b0;
        tmem_dat_o = 'b0;
        tmem_we_o  = 'b0;

        if (fu_i.ena) begin
            tmem_cyc_o = 1'b1;
            tmem_stb_o = 1'b1;
            tmem_adr_o = TADR_WIDTH'(mem_adr / GRANULARITY);

            case (fu_i.op)
                MTAG_OP_TADR: begin
                    tmem_dat_o = r_tag;
                    tmem_sel_o = '1;
                    tmem_we_o  = 'b1;
                end
                MTAG_OP_TADRE: begin
                    /* set tag in tag memory */
                    tmem_dat_o = enc_tag;
                    tmem_sel_o = '1;
                    tmem_we_o  = 'b1;
                end
                default: begin
                    /* unknown opcode */
                    err = 'b1;
                end
            endcase
        end
    end

    // output
    always_comb begin
        fu_o = funit_out_default();

        if (fu_i.ena) begin
            fu_o.rdy = 1'b1;
            fu_o.err = err;
        end
    end

endmodule
