// SPDX-License-Identifier: BSD-3-clause
/*
 * Copyright (C) Jörn Hoffmann, 2023
 *
 * Project  : SEC-V
 * Author   : J. Hoffmann <joern@bitaggregat.de>
 * Purpose  : Arithmetic-logic unit for the SEC-V processor.
 *
 * Opcodes
 *  - 64-Bit: ADD, SUB, SLL, SRL, SRA, SLT, SLTU, AND, OR, XOR
 *  - 32-Bit: ADDW, SUBW, SLLW, SRLW, SRAW
 *
 * Todo
 *  [ ] Add unit tests
 *  [ ] Add formal verification
 *
 * History
 *  v1.0    - Initial version
 */

`include "secv_pkg.svh"
import secv_pkg::*;

module alu #(
    parameter int XLEN = secv_pkg::XLEN
) (
    input  funit_in_t  fu_i,
    output funit_out_t fu_o
);

    logic [XLEN-1 : 0] res;
    logic err;

    alu_core #(
        .XLEN (XLEN)
    ) alu0 (
        .op_i   (fu_i.op),
        .a_i    (fu_i.src1),
        .b_i    (fu_i.src2),
        .res_o  (res)
    );

    // Output
    always_comb begin
        fu_o = funit_out_default();

        // Assign output, if unit is enabled and no error occured.
        // Unit is ready as soon as enabled.
        if (fu_i.ena) begin
            fu_o.rdy    = 1'b1;
            fu_o.err    = err;
            fu_o.res    = res;
            fu_o.res_wb = !err;
        end
    end
endmodule
